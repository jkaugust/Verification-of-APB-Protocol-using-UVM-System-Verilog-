module apb_slave (clk,rst,addr_in,wr,
