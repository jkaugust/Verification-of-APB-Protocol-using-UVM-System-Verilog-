module apb_master (clk,rst,addr_in,wr_in,ready,sel,
        data_in,sel_port,en,wr_out,addr_out,data_out);
  input clk;
  input rst;
  input [7:0] addr_in;
  input wr_in; //write when 1 and read when 0
  input ready;
  input sel;
  input [31:0] data_in;
  output reg [1:0] sel_port;
  output reg en;
  output reg wr_out;
  output reg [7:0] addr_out;
  output reg [31:0] data_out;
  
  reg [1:0] state;
 
  localparam [1:0]  IDLE    = 2'b00,
                    SETUP   = 2'b01,
                    ACCESS  = 2'b10,
                    WAIT    = 2'b11;
                    
                    
  always @(posedge clk)
    begin
      if (rst == 0) 
        begin 
          state    <= IDLE;
          addr_out <= 8'b0;
          data_out <= 32'b0;
          sel_port <= 2'b0;
          en       <= 0;
          wr_out   <= 0;   
        end
    else
      begin
        case (state)
          IDLE: begin
            addr_out   <= 8'b0;
            data_out   <= 32'b0;
            sel_port   <= 2'b0;
            en         <= 0;
            wr_out     <= 0;
            if (sel == 1) begin
              state  <= SETUP;
              end
              else begin
                state <= IDLE;
              end
            end
            
            SETUP: begin           
              sel_port   <= {>>{addr_in[7],addr_in[6]}};;
              en         <= 1;
              if (sel == 1) begin
                 state  <= ACCESS;
                end
                  else begin
                  state <= SETUP;
                end
              end
                
            ACCESS: begin
              if (ready == 1)
                begin
                  wr_out <= wr_in;
                  addr_out <= addr_in;
                  data_out <= data_in;
                  state <= WAIT;
                end
                  else begin
                  state <= ACCESS;
                end
              end
              
            
            WAIT: begin
                 en <= 0;
                if (sel == 1)
                  begin
                    if (ready == 0)
                      begin
                      state <= SETUP;
                      addr_out   <= 8'b0;
                      data_out   <= 32'b0;
                      sel_port   <= 2'b0;
                      wr_out     <= 0;
                     end
                   else
                     begin
                     state <= WAIT;
                    end
                  end
                else 
                  begin                     
                    state <= IDLE;
                  end
                end
                
              default: begin
                state <= IDLE;
              end
            endcase
          end
        end
 
  
endmodule
      




